 module Fetch(
	input CLK,
	output reg[19:0] INS
	);


