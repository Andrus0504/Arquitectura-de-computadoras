module module_and(
	input a,
	input b,
	output s);
assign s = a & b;
endmodule